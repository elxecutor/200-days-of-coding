Investigating Op-Amp Slew-Rate Limiting

* op-amp subcircuit
.subckt large_signal_opamp 1 2 3 6 4
* connections: | | | | |
* output | | \ /
* +ve input | |
* -ve input |
* current monitor of 1st stage
Iopen1 2 0 0A ; redundant connection made at +ve input terminal
Iopen2 3 0 0A ; redundant connection made at -ve input terminal
R 4 0 2.5Meg
C 4 5 30p
Ginput 6 0 Table {V(2)-V(3)} = (-0.1V,-19uA) (0.1V,19uA)
Emiddle 5 0 4 0 -529
Eoutput 1 0 Table {V(5)} = (-10V,-10V) (10V,10V)
.ends large_signal_opamp

** Main Circuit **
* signal source
Vi 2 0 PWL (0,0V 1us,0V 1.01us,1mV 1s,1mV )
Xopamp 1 2 1 4 5 large_signal_opamp
Vmonitor 4 5 0

** Analysis Requests **
.TRAN 10ns 5us 0s 10ns
** Output Requests **
.PLOT TRAN V(2) V(1) I(Vmonitor)
.probe
.end
