Investigating The Sensitivity Of the Emitter Current To Amplifier Components

** Circuit Description **
* power supply
Vcc 1 0 DC +12V
* amplifier circuit
Q1 2 3 4 Q2N2222A
Rc 1 2 4k
R1 1 3 80k
R2 3 0 40k
Re 4 5 3.3k
Vemitter 5 0 0
* transistor model statement for the 2N2222A
.model Q2N2222A NPN (Is=14.34f Xti=3 Eg=1.11 Vaf=74.03 Bf=255.9 Ne=1.307
+                    Ise=14.34f Ikf=.2847 Xtb=1.5 Br=6.092 Nc=2 Isc=0 Ikr=0 Rc=1
+                    Cjc=7.306p Mjc=.3416 Vjc=.75 Fc=.5 Cje=22.01p Mje=.377 Vje=.75
+                    Tr=46.91n Tf=411.1p Itf=.6 Vtf=1.7 Xtf=3 Rb=10)
** Analysis Requests **
.op
** Output Requests **
* none required
.end
