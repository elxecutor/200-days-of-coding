** Circuit Description **

* signal source
Vi 3 0 DC 1v
* inverting amplifier circuit description
R1 3 2 1k
R2 2 1 10k
Eopamp 1 0 0 2 1e6

** Analysis Requests **
.TF V(1) Vi

** Output Requests **
* none required

.end
